module partial_product_28bit
(
	output [27:0]out,
	input  [27:0]x,
	input   y
);
	and (out[0], x[0], y);
	and (out[1], x[1], y);
	and (out[2], x[2], y);
	and (out[3], x[3], y);
	and (out[4], x[4], y);
	and (out[5], x[5], y);
	and (out[6], x[6], y);
	and (out[7], x[7], y);
	and (out[8], x[8], y);
	and (out[9], x[9], y);
	and (out[10], x[10], y);
	and (out[11], x[11], y);
	and (out[12], x[12], y);
	and (out[13], x[13], y);
	and (out[14], x[14], y);
	and (out[15], x[15], y);
	and (out[16], x[16], y);
	and (out[17], x[17], y);
	and (out[18], x[18], y);
	and (out[19], x[19], y);
	and (out[20], x[20], y);
	and (out[21], x[21], y);
	and (out[22], x[22], y);
	and (out[23], x[23], y);
	and (out[24], x[24], y);
	and (out[25], x[25], y);
	and (out[26], x[26], y);
	and (out[27], x[27], y);


endmodule
