module Butterfly(
    output [24-1:0] C1, C2,
    input [24-1:0] A, B
);

    assign C1[23:12] = ({A[23], A[23:12]} + {B[23], B[23:12]}) >> 1;
    assign C1[11:0] = ({A[11], A[11:0]} + {B[11], B[11:0]}) >> 1;
    assign C2[23:12] = ({A[23], A[23:12]} - {B[23], B[23:12]}) >> 1;
    assign C2[11:0] = ({A[11], A[11:0]} - {B[11], B[11:0]}) >> 1;

endmodule
